--============================================================================--
-- Design unit  : rom_data
--
-- File name    : Rom_256n08.vhd
--
-- Purpose      : data for the ROM
--
-- Note         :
--
-- Library      : shyloc_utils
--
-- Author       : Rui Yin
--
-- Instantiates : 
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

package ROM_Package is
	
	constant width	: integer := 32;
        constant depth : integer:= 128;
	constant addr : integer := 8;
    type ROM_ARRAY is array (0 to depth-1) of STD_LOGIC_VECTOR(width-1 downto 0);
    constant ROM_CONTENT: ROM_ARRAY := (
    0 => X"FF7FFEFF",
    1 => X"FF7FFFFF",
    2 => X"FF7F0000",
    3 => X"0080FFFF",
    4 => X"00800100",
    5 => X"00800000",
    6 => X"FF7FFDFF",
    7 => X"0000FFFF",
    8 => X"00000060",
    9 => X"00200020",
    10 => X"00500010",
    11 => X"00100040",
    12 => X"00000000",
    13 => X"00600020",
    14 => X"00200050",
    15 => X"00100010",
    16 => X"00000020",
    17 => X"00300040",
    18 => X"00500060",
    19 => X"00700080",
    20 => X"00900070",
    21 => X"00600050",
    22 => X"00400030",
    23 => X"00200010",
    24 => X"00200020",
    25 => X"00300040",
    26 => X"00500060",
    27 => X"00700080",
    28 => X"00900070",
    29 => X"00600050",
    30 => X"00400030",
    31 => X"00200020",
    32 => X"00100010",
    33 => X"00180020",
    34 => X"00280030",
    35 => X"00380040",
    36 => X"00480038",
    37 => X"00300028",
    38 => X"00200018",
    39 => X"00100010",
    40 => X"00080008",
    41 => X"000C0010",
    42 => X"00140018",
    43 => X"001C0020",
    44 => X"0024001C",
    45 => X"00180014",
    46 => X"0010000C",
    47 => X"00080008",
    48 => X"00040004",
    49 => X"00060008",
    50 => X"000A000C",
    51 => X"000E0010",
    52 => X"0012000E",
    53 => X"000C000A",
    54 => X"00080006",
    55 => X"00040004",
    56 => X"00020002",
    57 => X"00030004",
    58 => X"00050006",
    59 => X"00070008",
    60 => X"00090007",
    61 => X"00060005",
    62 => X"00040003",
    63 => X"00020002",
    64 => X"00010001",
    65 => X"80010002",
    66 => X"80020003",
    67 => X"80030004",
    68 => X"80048003",
    69 => X"00038002",
    70 => X"00028001",
    71 => X"00010001",
    72 => X"80008000",
    73 => X"C0000001",
    74 => X"40018001",
    75 => X"C0010002",
    76 => X"4002C001",
    77 => X"80014001",
    78 => X"0001C000",
    79 => X"80008000",
    80 => X"40004000",
    81 => X"60008000",
    82 => X"A000C000",
    83 => X"E0000001",
    84 => X"2001E000",
    85 => X"C000A000",
    86 => X"80006000",
    87 => X"40004000",
    88 => X"20002000",
    89 => X"30004000",
    90 => X"50006000",
    91 => X"70008000",
    92 => X"90007000",
    93 => X"60005000",
    94 => X"40003000",
    95 => X"20002000",
    96 => X"10001000",
    97 => X"18002000",
    98 => X"28003000",
    99 => X"38004000",
    100 => X"48003800",
    101 => X"30002800",
    102 => X"20001800",
    103 => X"10001000",
    104 => X"08000800",
    105 => X"0C001000",
    106 => X"14001800",
    107 => X"1C002000",
    108 => X"24001C00",
    109 => X"18001400",
    110 => X"10000C00",
    111 => X"08000800",
    112 => X"04000400",
    113 => X"06000800",
    114 => X"0A000C00",
    115 => X"0E001000",
    116 => X"12000E00",
    117 => X"0C000A00",
    118 => X"08000600",
    119 => X"04000400",
    120 => X"02000200",
    121 => X"03000400",
    122 => X"05000600",
    123 => X"07000800",
    124 => X"09000700",
    125 => X"06000500",
    126 => X"04000300",
    127 => X"02000200",
	others => (others => '0'));
end ROM_Package;
